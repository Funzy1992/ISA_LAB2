//`timescale 1ns

module tb_fir ();

   wire CLK_i;
   wire RST_n_i;
   wire [7:0] DIN_0i;
   wire [7:0] DIN_1i;
   wire [7:0] DIN_2i;
   wire [7:0] DOUT_0i;
   wire [7:0] DOUT_1i;
   wire [7:0] DOUT_2i;
   wire VIN_i;
   wire signed [7:0] H0_i;
   wire signed [7:0] H1_i;
   wire signed [7:0] H2_i;
   wire signed [7:0] H3_i;
   wire signed [7:0] H4_i;
   wire signed [7:0] H5_i;
   wire signed [7:0] H6_i;
   wire signed [7:0] H7_i;
   wire signed [7:0] H8_i;
   wire signed [7:0] H9_i;
   wire signed [7:0] H10_i;
   wire [7:0] DOUT_i;
   wire VOUT_i;
   wire END_SIM_i;

   clk_gen CG(.END_SIM(END_SIM_i),
  	      .CLK(CLK_i),
	      .RST_n(RST_n_i));

   data_maker SM(.CLK(CLK_i),
	         .RST_n(RST_n_i),
			 .VOUT(VIN_i),
			 .DOUT_0(DIN_0i),
			 .DOUT_1(DIN_1i),
			 .DOUT_2(DIN_2i),
			 .H0(H0_i),
			 .H1(H1_i),
			 .H2(H2_i),
			 .H3(H3_i),
			 .H4(H4_i),
			 .H5(H5_i),
			 .H6(H6_i),
			 .H7(H7_i),
			 .H8(H8_i),
			 .H9(H9_i),
			 .H10(H10_i),
			 .END_SIM(END_SIM_i));

   Unfolded_FIR UUT(.CLK(CLK_i),
	     .RESET(RST_n_i),			//reset=rst_n
		 .VIN(VIN_i),
	     .B0(H0_i),
	     .B1(H1_i),
	     .B2(H2_i),
	     .B3(H3_i),
		 .B4(H4_i),
		 .B5(H5_i),
		 .B6(H6_i),
		 .B7(H7_i),
		 .B8(H8_i),
		 .B9(H9_i),
		 .B10(H10_i),
		 .DIN_0(DIN_0i),
		 .DIN_1(DIN_1i),
		 .DIN_2(DIN_2i),
		 .DOUT_0(DOUT_0i),
		 .DOUT_1(DOUT_1i),
		 .DOUT_2(DOUT_2i),		 
		 .VOUT(VOUT_i));

   data_sink DS(.CLK(CLK_i),
		.RST_n(RST_n_i),
		.VIN(VOUT_i),
		.DIN_0(DOUT_0i),
		.DIN_1(DOUT_1i),
		.DIN_2(DOUT_2i));   

endmodule

		   